class transaction;
rand bit [7:0] din;
rand bit [7:0] addr;
bit wr;
bit [7:0] dout;
endclass
