interface counter_intf();
logic clk, rst, wr;
logic [7:0] din, addr;
logic [7:0] dout;
endinterface
 
